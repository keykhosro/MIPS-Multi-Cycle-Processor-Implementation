library verilog;
use verilog.vl_types.all;
entity multiplier is
    port(
        clk             : in     vl_logic;
        start           : in     vl_logic;
        A               : in     vl_logic_vector(31 downto 0);
        B               : in     vl_logic_vector(31 downto 0);
        Product         : out    vl_logic_vector(63 downto 0);
        ready           : out    vl_logic
    );
end multiplier;
